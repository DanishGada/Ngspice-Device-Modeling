su
.subckt nandcmos a b y
vdd 1 0 dc 5v
m1 1 a y 1 mos1 l=10u w=100u
m2 1 b y 1 mos1 l=10u w=100u
m3 y a 2 0 mos2 l=10u w=100u
m4 2 b 0 0 mos2 l=10u w=100u
.model mos1 pmos vto=1.5v kp=200u
.model mos2 nmos vto=1.5v kp=200u
.ends

.subckt notcmos a y
vdd 1 0 dc 5v
m1 1 a y 1 mos1 l=10u w=100u
m2 y a 0 0 mos2 l=10u w=100u
.model mos1 pmos vt0=1.5v kp=200u
.model mos2 nmos vt0=1.5v kp=200u
.ends
.subckt kuchtohincmos a b y
vdd 1 0 dc 5v
m1 1 a y 1 mos1 l=10u w=100u
m2 y a b b mos2 l=10u w=100u
.model mos1 pmos vt0=1.5v kp=200u
.model mos2 nmos vt0=1.5v kp=200u
.ends

Va a 0 pulse(0 5 0 0 0 10s 20s)
Vb b 0 pulse(0 5 0 0 0 20s 40s)
X1 b y notcmos
X2 a y z2 kuchtohincmos
X3 a b z1 nandcmos

.control
tran 0.1s 40s
plot v(a) v(b)+6 v(z1)+12 v(z2)+24
.endc
.end